module chacha20

